*** Input filter (real op-amp) ***

* Input audio source
* See https://en.wikipedia.org/wiki/Line_level
vin inp inn 0 dc 1.414 ac

.include analog_input_buffer.cir
x2a 2 4 V12+ V12- 5 OPA1622
x2b 3 7 V12+ V12- 8 OPA1622
.include OPA1622.txt

* let's analyze the frequency response
.ac dec 100 1 20Meg

.end
