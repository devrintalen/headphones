CS5381 input filter (real op-amp and real caps)

* Capacitor selections
*
* c11/12 : C2012X7R1A106K125AC
* c13/14 : C2012C0G2W471J060AA
* c15    : C2012X7R1H104K085AA
* c16    : C2012C0G1H272J060AA
* 

vin inp inn 0 dc 1.414 ac sin(0 1.414 1K)
v12p V12+ 0 dc 12V trnoise(10m 10u 0 0)
v12n V12- 0 dc -12V trnoise(10m 10u 0 0)
vqst VQ   0 dc 2.5V trnoise(10m 10u 0 0)

r5 inp 0 100Kohm
r7 2 VQ 10Kohm
r99 inn 0 0ohm
r6 inn 0 100Kohm
r8 3 VQ 10Kohm
r11 5 6 91ohm
r9  4 6 634ohm
r13 6 ainp 200ohm
r12 8 9 91ohm
r10 7 9 634ohm
r14 9 ainn 200ohm
r15 ainp ainn 200ohm

x11 2    inp  C2012X7R1A106K125AC_p
x12 3    inn  C2012X7R1A106K125AC_p
x13 4    5    C2012C0G2W471J060AA_p
x14 7    8    C2012C0G2W471J060AA_p
x15 VQ   0    C2012X7R1H104K085AA_p
x16 ainp ainn C2012C0G1H272J060AA_p

.include C2012C0G1H272J060AA_p.mod
.include C2012C0G2W471J060AA_p.mod
.include C2012X7R1H104K085AA_p.mod
.include C2012X7R1A106K125AC_p.mod

x2a 2 4 V12+ V12- 5 OPA1622
x2b 3 7 V12+ V12- 8 OPA1622

.func LIMIT(x,a,b) {min(max(x, a), b)}
.func PWR(x,a) {abs(x) ** a}
.func PWRS(x,a) {sgn(x) * PWR(x,a)}
.func stp(x) {u(x)}
.include OPA1622.txt

.control
set noaskquit
ac dec 100 1 20Meg
wrdata adc_precise_ac db( v(ainp,ainn) / v(inp,inn) )
tran 10u 20m 0m 10u
fourier 1K v(ainp,ainn)
wrdata adc_precise_tran v(ainp,ainn) v(inp,inn)
let vout = v(ainp,ainn)
spec 20 20K 50 vout
wrdata adc_precise_spec mag(vout)
quit
.endc

.end
