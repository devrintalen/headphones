CS5381 input filter (ideal)

vin inp inn 0 dc 1.414 ac sin(0 1.414 1K)
v12p V12+ 0 dc 12V
v12n V12- 0 dc -12V
vqst VQ   0 dc 2.5V

r5 inp 0 100Kohm
c11 2 inp 10uF
r7 2 VQ 10Kohm
c15 VQ 0 0.1uF
r99 inn 0 0ohm
r6 inn 0 100Kohm
c12 3 inn 10uF
r8 3 VQ 10Kohm
c13 4 5 470pF
r11 5 6 91ohm
r9  4 6 634ohm
r13 6 ainp 200ohm
C14 7 8 470pF
r12 8 9 91ohm
r10 7 9 634ohm
r14 9 ainn 200ohm
r15 ainp ainn 200ohm
c16 ainp ainn 2700pF

x2a 2 4 V12+ V12- 5 LM741/NS
x2b 3 7 V12+ V12- 8 LM741/NS
.include LM741.MOD

.control
set noaskquit
ac dec 100 1 20Meg
wrdata adc_ideal_ac db( v(ainp,ainn) / v(inp,inn) )
tran 10u 20m 0m 10u
fourier 1K v(ainp,ainn)
wrdata adc_ideal_tran v(ainp,ainn) v(inp,inn)
let vout = v(ainp,ainn)
spec 20 20K 50 vout
wrdata adc_ideal_spec mag(vout)
quit
.endc

.end
